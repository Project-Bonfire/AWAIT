--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated Please do not change!
-- Here are the parameters:
-- 	 network size x:4
-- 	 network size y:4
-- 	 data width:32-- 	 traffic pattern:------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.TB_Package.all;
use work.component_pack.all;

USE ieee.numeric_std.ALL; 
use IEEE.math_real."ceil";
use IEEE.math_real."log2";

entity tb_router is
    --Pass the filenames to write to for the sent and received file.
	--generic (sent_file,recv_file : string);
end tb_router; 

architecture behavior of tb_router is

    -- generating bulk signals...

    --define the signals of the router
	signal RX_L_5, TX_L_5, 
           RX_N_5, RX_E_5, RX_W_5, RX_S_5,	
		   TX_N_5, TX_E_5, TX_W_5, TX_S_5:  std_logic_vector (31 downto 0);

	signal credit_in_N_5, credit_in_E_5, credit_in_W_5, credit_in_S_5, credit_in_L_5, 
           valid_in_N_5, valid_in_E_5, valid_in_W_5, valid_in_S_5, valid_in_L_5,
		   valid_out_N_5, valid_out_E_5, valid_out_W_5, valid_out_S_5, valid_out_L_5,
		   credit_out_N_5, credit_out_E_5, credit_out_W_5, credit_out_S_5, credit_out_L_5: std_logic;

    signal Faulty_in_N_5, Faulty_in_E_5, Faulty_in_W_5, Faulty_in_S_5: std_logic := '0';
    signal Faulty_out_N_5, Faulty_out_E_5, Faulty_out_W_5, Faulty_out_S_5: std_logic;

	signal credit_counter_out_5:  std_logic_vector (1 downto 0);
	signal credit_counter_out_1:  std_logic_vector (1 downto 0);
	signal credit_counter_out_4:  std_logic_vector (1 downto 0);
	signal credit_counter_out_6:  std_logic_vector (1 downto 0);
	signal credit_counter_out_9:  std_logic_vector (1 downto 0);

	--------------
    signal Rxy_reconf_PE_5: std_logic_vector (7 downto 0) := "00111100";
    signal Cx_reconf_PE_5:  std_logic_vector (3 downto 0) := "1111";
	signal Reconfig_command_5: std_logic := '0';

    signal link_faults_5: std_logic_vector (4 downto  0);
    signal turn_faults_5: std_logic_vector (19 downto 0);

    signal link_faults_async_5: std_logic_vector (4 downto  0);
    signal turn_faults_async_5: std_logic_vector (19 downto 0);

	--------------
	constant clk_period : time := 10 ns;
	signal reset, not_reset, clk: std_logic :='0';

begin

   clk_process :process
   begin
        clk <= '0';
        wait for clk_period/2;   
        clk <= '1';
        wait for clk_period/2; 
   end process;

reset <= '1' after 1 ns;


-- instantiating the router

R_5: router_credit_based_PD_C_SHMU_with_checkers
generic map (DATA_WIDTH => 32, current_address => 5, Rxy_rst => 60, Cx_rst => 15, healthy_counter_threshold => 15, faulty_counter_threshold => 4, counter_depth => 4, NoC_size => 4)
PORT MAP (  reset, clk, 

        	RX_N => RX_N_5, RX_E => RX_E_5, RX_W => RX_W_5, RX_S => RX_S_5, RX_L => RX_L_5,
        	credit_in_N => credit_in_N_5, credit_in_E => credit_in_E_5, credit_in_W => credit_in_W_5, credit_in_S => credit_in_S_5, credit_in_L => credit_in_L_5,
        	valid_in_N => valid_in_N_5, valid_in_E => valid_in_E_5, valid_in_W => valid_in_W_5, valid_in_S => valid_in_S_5, valid_in_L => valid_in_L_5,
        	valid_out_N => valid_out_N_5, valid_out_E => valid_out_E_5, valid_out_W => valid_out_W_5, valid_out_S => valid_out_S_5, valid_out_L => valid_out_L_5,
            credit_out_N => credit_out_N_5, credit_out_E => credit_out_E_5, credit_out_W => credit_out_W_5, credit_out_S => credit_out_S_5, credit_out_L => credit_out_L_5,
            TX_N => TX_N_5, TX_E => TX_E_5, TX_W => TX_W_5, TX_S => TX_S_5, TX_L => TX_L_5,

            Faulty_N_in => Faulty_in_N_5, Faulty_E_in => Faulty_in_E_5, Faulty_W_in => Faulty_in_W_5, Faulty_S_in => Faulty_in_S_5,  
            Faulty_N_out => Faulty_out_N_5, Faulty_E_out => Faulty_out_E_5, Faulty_W_out => Faulty_out_W_5, Faulty_S_out => Faulty_out_S_5, 

            link_faults => link_faults_5, 
            turn_faults => turn_faults_5, 

            Rxy_reconf_PE => Rxy_reconf_PE_5, 
            Cx_reconf_PE => Cx_reconf_PE_5, 
            Reconfig_command => Reconfig_command_5, 

            link_faults_async => link_faults_async_5, 
            turn_faults_async => turn_faults_async_5
         ); 

not_reset <= not reset; 

-- connecting the packet generators
 
--set up traffic generators
credit_counter_control(clk, credit_out_L_5, valid_in_L_5, credit_counter_out_5);
gen_random_packet("sent.txt",4, 50, 5, 23, 8, 8, 10000 ns, clk, credit_counter_out_5, valid_in_L_5, RX_L_5);

credit_counter_control(clk, credit_out_N_5, valid_in_N_5, credit_counter_out_1);
gen_random_packet("sent.txt",4, 50, 1, 23, 8, 8, 10000 ns, clk, credit_counter_out_1, valid_in_N_5, RX_N_5);

credit_counter_control(clk, credit_out_E_5, valid_in_E_5, credit_counter_out_6);
gen_random_packet("sent.txt",4, 50, 6, 23, 8, 8, 10000 ns, clk, credit_counter_out_6, valid_in_E_5, RX_E_5);

credit_counter_control(clk, credit_out_S_5, valid_in_S_5, credit_counter_out_9);
gen_random_packet("sent.txt",4, 50, 9, 23, 8, 8, 10000 ns, clk, credit_counter_out_9, valid_in_S_5, RX_S_5);

credit_counter_control(clk, credit_out_W_5, valid_in_W_5, credit_counter_out_4);
gen_random_packet("sent.txt",4, 50, 4, 23, 8, 8, 10000 ns, clk, credit_counter_out_4, valid_in_W_5, RX_W_5);



-- connecting the packet receivers
get_packet("received.txt",32, 5, 1, clk, credit_in_N_5, valid_out_N_5, TX_N_5);
get_packet("received.txt",32, 5, 6, clk, credit_in_E_5, valid_out_E_5, TX_E_5);
get_packet("received.txt",32, 5, 9, clk, credit_in_S_5, valid_out_S_5, TX_S_5);
get_packet("received.txt",32, 5, 4, clk, credit_in_W_5, valid_out_W_5, TX_W_5);
get_packet("received.txt",32, 5, 5, clk, credit_in_L_5, valid_out_L_5, TX_L_5);


end;
