--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated Please do not change!
-- Here are the parameters:
-- 	 network size x:4
-- 	 network size y:4
-- 	 data width:32-- 	 traffic pattern:------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.TB_Package.all;

--use work.router_pack.all;

USE ieee.numeric_std.ALL; 
use IEEE.math_real."ceil";
use IEEE.math_real."log2";

entity tb_network_4x4 is
end tb_network_4x4; 


architecture behavior of tb_network_4x4 is

-- Declaring network component
component network_4x4 is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic; 
	clk: in  std_logic; 
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_0, valid_out_L_0: out std_logic;
	credit_in_L_0, valid_in_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_1, valid_out_L_1: out std_logic;
	credit_in_L_1, valid_in_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_2, valid_out_L_2: out std_logic;
	credit_in_L_2, valid_in_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_3, valid_out_L_3: out std_logic;
	credit_in_L_3, valid_in_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_4: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_4, valid_out_L_4: out std_logic;
	credit_in_L_4, valid_in_L_4: in std_logic;
	TX_L_4: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_5: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_5, valid_out_L_5: out std_logic;
	credit_in_L_5, valid_in_L_5: in std_logic;
	TX_L_5: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_6: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_6, valid_out_L_6: out std_logic;
	credit_in_L_6, valid_in_L_6: in std_logic;
	TX_L_6: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_7: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_7, valid_out_L_7: out std_logic;
	credit_in_L_7, valid_in_L_7: in std_logic;
	TX_L_7: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_8: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_8, valid_out_L_8: out std_logic;
	credit_in_L_8, valid_in_L_8: in std_logic;
	TX_L_8: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_9: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_9, valid_out_L_9: out std_logic;
	credit_in_L_9, valid_in_L_9: in std_logic;
	TX_L_9: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_10: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_10, valid_out_L_10: out std_logic;
	credit_in_L_10, valid_in_L_10: in std_logic;
	TX_L_10: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_11: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_11, valid_out_L_11: out std_logic;
	credit_in_L_11, valid_in_L_11: in std_logic;
	TX_L_11: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_12: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_12, valid_out_L_12: out std_logic;
	credit_in_L_12, valid_in_L_12: in std_logic;
	TX_L_12: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_13: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_13, valid_out_L_13: out std_logic;
	credit_in_L_13, valid_in_L_13: in std_logic;
	TX_L_13: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_14: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_14, valid_out_L_14: out std_logic;
	credit_in_L_14, valid_in_L_14: in std_logic;
	TX_L_14: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_15: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_15, valid_out_L_15: out std_logic;
	credit_in_L_15, valid_in_L_15: in std_logic;
	TX_L_15: out std_logic_vector (DATA_WIDTH-1 downto 0); 

	--------------
    link_faults_0: out std_logic_vector(4 downto 0);
    turn_faults_0: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_0: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_0: in  std_logic_vector(3 downto 0);
    Reconfig_command_0 : in std_logic;
    link_faults_async_0: out std_logic_vector(4 downto 0);
    turn_faults_async_0: out std_logic_vector(19 downto 0);

	--------------
    link_faults_1: out std_logic_vector(4 downto 0);
    turn_faults_1: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_1: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_1: in  std_logic_vector(3 downto 0);
    Reconfig_command_1 : in std_logic;
    link_faults_async_1: out std_logic_vector(4 downto 0);
    turn_faults_async_1: out std_logic_vector(19 downto 0);

	--------------
    link_faults_2: out std_logic_vector(4 downto 0);
    turn_faults_2: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_2: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_2: in  std_logic_vector(3 downto 0);
    Reconfig_command_2 : in std_logic;
    link_faults_async_2: out std_logic_vector(4 downto 0);
    turn_faults_async_2: out std_logic_vector(19 downto 0);

	--------------
    link_faults_3: out std_logic_vector(4 downto 0);
    turn_faults_3: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_3: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_3: in  std_logic_vector(3 downto 0);
    Reconfig_command_3 : in std_logic;
    link_faults_async_3: out std_logic_vector(4 downto 0);
    turn_faults_async_3: out std_logic_vector(19 downto 0);

	--------------
    link_faults_4: out std_logic_vector(4 downto 0);
    turn_faults_4: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_4: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_4: in  std_logic_vector(3 downto 0);
    Reconfig_command_4 : in std_logic;
    link_faults_async_4: out std_logic_vector(4 downto 0);
    turn_faults_async_4: out std_logic_vector(19 downto 0);

	--------------
    link_faults_5: out std_logic_vector(4 downto 0);
    turn_faults_5: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_5: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_5: in  std_logic_vector(3 downto 0);
    Reconfig_command_5 : in std_logic;
    link_faults_async_5: out std_logic_vector(4 downto 0);
    turn_faults_async_5: out std_logic_vector(19 downto 0);

	--------------
    link_faults_6: out std_logic_vector(4 downto 0);
    turn_faults_6: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_6: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_6: in  std_logic_vector(3 downto 0);
    Reconfig_command_6 : in std_logic;
    link_faults_async_6: out std_logic_vector(4 downto 0);
    turn_faults_async_6: out std_logic_vector(19 downto 0);

	--------------
    link_faults_7: out std_logic_vector(4 downto 0);
    turn_faults_7: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_7: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_7: in  std_logic_vector(3 downto 0);
    Reconfig_command_7 : in std_logic;
    link_faults_async_7: out std_logic_vector(4 downto 0);
    turn_faults_async_7: out std_logic_vector(19 downto 0);

	--------------
    link_faults_8: out std_logic_vector(4 downto 0);
    turn_faults_8: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_8: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_8: in  std_logic_vector(3 downto 0);
    Reconfig_command_8 : in std_logic;
    link_faults_async_8: out std_logic_vector(4 downto 0);
    turn_faults_async_8: out std_logic_vector(19 downto 0);

	--------------
    link_faults_9: out std_logic_vector(4 downto 0);
    turn_faults_9: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_9: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_9: in  std_logic_vector(3 downto 0);
    Reconfig_command_9 : in std_logic;
    link_faults_async_9: out std_logic_vector(4 downto 0);
    turn_faults_async_9: out std_logic_vector(19 downto 0);

	--------------
    link_faults_10: out std_logic_vector(4 downto 0);
    turn_faults_10: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_10: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_10: in  std_logic_vector(3 downto 0);
    Reconfig_command_10 : in std_logic;
    link_faults_async_10: out std_logic_vector(4 downto 0);
    turn_faults_async_10: out std_logic_vector(19 downto 0);

	--------------
    link_faults_11: out std_logic_vector(4 downto 0);
    turn_faults_11: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_11: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_11: in  std_logic_vector(3 downto 0);
    Reconfig_command_11 : in std_logic;
    link_faults_async_11: out std_logic_vector(4 downto 0);
    turn_faults_async_11: out std_logic_vector(19 downto 0);

	--------------
    link_faults_12: out std_logic_vector(4 downto 0);
    turn_faults_12: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_12: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_12: in  std_logic_vector(3 downto 0);
    Reconfig_command_12 : in std_logic;
    link_faults_async_12: out std_logic_vector(4 downto 0);
    turn_faults_async_12: out std_logic_vector(19 downto 0);

	--------------
    link_faults_13: out std_logic_vector(4 downto 0);
    turn_faults_13: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_13: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_13: in  std_logic_vector(3 downto 0);
    Reconfig_command_13 : in std_logic;
    link_faults_async_13: out std_logic_vector(4 downto 0);
    turn_faults_async_13: out std_logic_vector(19 downto 0);

	--------------
    link_faults_14: out std_logic_vector(4 downto 0);
    turn_faults_14: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_14: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_14: in  std_logic_vector(3 downto 0);
    Reconfig_command_14 : in std_logic;
    link_faults_async_14: out std_logic_vector(4 downto 0);
    turn_faults_async_14: out std_logic_vector(19 downto 0);

	--------------
    link_faults_15: out std_logic_vector(4 downto 0);
    turn_faults_15: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_15: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_15: in  std_logic_vector(3 downto 0);
    Reconfig_command_15 : in std_logic;
    link_faults_async_15: out std_logic_vector(4 downto 0);
    turn_faults_async_15: out std_logic_vector(19 downto 0);

    -- for bubbles
    --------------
    hold_in_N_0, hold_in_E_0, hold_in_S_0, hold_in_W_0, hold_in_L_0: in std_logic;
    hold_out_N_0, hold_out_E_0, hold_out_S_0, hold_out_W_0, hold_out_L_0: out std_logic;

	--------------
    hold_in_N_1, hold_in_E_1, hold_in_S_1, hold_in_W_1, hold_in_L_1: in std_logic;
    hold_out_N_1, hold_out_E_1, hold_out_S_1, hold_out_W_1, hold_out_L_1: out std_logic;

	--------------
    hold_in_N_2, hold_in_E_2, hold_in_S_2, hold_in_W_2, hold_in_L_2: in std_logic;
    hold_out_N_2, hold_out_E_2, hold_out_S_2, hold_out_W_2, hold_out_L_2: out std_logic;

	--------------
    hold_in_N_3, hold_in_E_3, hold_in_S_3, hold_in_W_3, hold_in_L_3: in std_logic;
    hold_out_N_3, hold_out_E_3, hold_out_S_3, hold_out_W_3, hold_out_L_3: out std_logic;

	--------------
    hold_in_N_4, hold_in_E_4, hold_in_S_4, hold_in_W_4, hold_in_L_4: in std_logic;
    hold_out_N_4, hold_out_E_4, hold_out_S_4, hold_out_W_4, hold_out_L_4: out std_logic;

	--------------
    hold_in_N_5, hold_in_E_5, hold_in_S_5, hold_in_W_5, hold_in_L_5: in std_logic;
    hold_out_N_5, hold_out_E_5, hold_out_S_5, hold_out_W_5, hold_out_L_5: out std_logic;

	--------------
    hold_in_N_6, hold_in_E_6, hold_in_S_6, hold_in_W_6, hold_in_L_6: in std_logic;
    hold_out_N_6, hold_out_E_6, hold_out_S_6, hold_out_W_6, hold_out_L_6: out std_logic;

	--------------
    hold_in_N_7, hold_in_E_7, hold_in_S_7, hold_in_W_7, hold_in_L_7: in std_logic;
    hold_out_N_7, hold_out_E_7, hold_out_S_7, hold_out_W_7, hold_out_L_7: out std_logic;

	--------------
    hold_in_N_8, hold_in_E_8, hold_in_S_8, hold_in_W_8, hold_in_L_8: in std_logic;
    hold_out_N_8, hold_out_E_8, hold_out_S_8, hold_out_W_8, hold_out_L_8: out std_logic;

	--------------
    hold_in_N_9, hold_in_E_9, hold_in_S_9, hold_in_W_9, hold_in_L_9: in std_logic;
    hold_out_N_9, hold_out_E_9, hold_out_S_9, hold_out_W_9, hold_out_L_9: out std_logic;

	--------------
    hold_in_N_10, hold_in_E_10, hold_in_S_10, hold_in_W_10, hold_in_L_10: in std_logic;
    hold_out_N_10, hold_out_E_10, hold_out_S_10, hold_out_W_10, hold_out_L_10: out std_logic;

	--------------
    hold_in_N_11, hold_in_E_11, hold_in_S_11, hold_in_W_11, hold_in_L_11: in std_logic;
    hold_out_N_11, hold_out_E_11, hold_out_S_11, hold_out_W_11, hold_out_L_11: out std_logic;

	--------------
    hold_in_N_12, hold_in_E_12, hold_in_S_12, hold_in_W_12, hold_in_L_12: in std_logic;
    hold_out_N_12, hold_out_E_12, hold_out_S_12, hold_out_W_12, hold_out_L_12: out std_logic;

	--------------
    hold_in_N_13, hold_in_E_13, hold_in_S_13, hold_in_W_13, hold_in_L_13: in std_logic;
    hold_out_N_13, hold_out_E_13, hold_out_S_13, hold_out_W_13, hold_out_L_13: out std_logic;

	--------------
    hold_in_N_14, hold_in_E_14, hold_in_S_14, hold_in_W_14, hold_in_L_14: in std_logic;
    hold_out_N_14, hold_out_E_14, hold_out_S_14, hold_out_W_14, hold_out_L_14: out std_logic;

	--------------
    hold_in_N_15, hold_in_E_15, hold_in_S_15, hold_in_W_15, hold_in_L_15: in std_logic;
    hold_out_N_15, hold_out_E_15, hold_out_S_15, hold_out_W_15, hold_out_L_15: out std_logic

   ); 

end component; 

-- generating bulk signals...
	signal RX_L_0, TX_L_0:  std_logic_vector (31 downto 0);
	signal credit_counter_out_0:  std_logic_vector (1 downto 0);
	signal credit_out_L_0, credit_in_L_0, valid_in_L_0, valid_out_L_0: std_logic;
	signal RX_L_1, TX_L_1:  std_logic_vector (31 downto 0);
	signal credit_counter_out_1:  std_logic_vector (1 downto 0);
	signal credit_out_L_1, credit_in_L_1, valid_in_L_1, valid_out_L_1: std_logic;
	signal RX_L_2, TX_L_2:  std_logic_vector (31 downto 0);
	signal credit_counter_out_2:  std_logic_vector (1 downto 0);
	signal credit_out_L_2, credit_in_L_2, valid_in_L_2, valid_out_L_2: std_logic;
	signal RX_L_3, TX_L_3:  std_logic_vector (31 downto 0);
	signal credit_counter_out_3:  std_logic_vector (1 downto 0);
	signal credit_out_L_3, credit_in_L_3, valid_in_L_3, valid_out_L_3: std_logic;
	signal RX_L_4, TX_L_4:  std_logic_vector (31 downto 0);
	signal credit_counter_out_4:  std_logic_vector (1 downto 0);
	signal credit_out_L_4, credit_in_L_4, valid_in_L_4, valid_out_L_4: std_logic;
	signal RX_L_5, TX_L_5:  std_logic_vector (31 downto 0);
	signal credit_counter_out_5:  std_logic_vector (1 downto 0);
	signal credit_out_L_5, credit_in_L_5, valid_in_L_5, valid_out_L_5: std_logic;
	signal RX_L_6, TX_L_6:  std_logic_vector (31 downto 0);
	signal credit_counter_out_6:  std_logic_vector (1 downto 0);
	signal credit_out_L_6, credit_in_L_6, valid_in_L_6, valid_out_L_6: std_logic;
	signal RX_L_7, TX_L_7:  std_logic_vector (31 downto 0);
	signal credit_counter_out_7:  std_logic_vector (1 downto 0);
	signal credit_out_L_7, credit_in_L_7, valid_in_L_7, valid_out_L_7: std_logic;
	signal RX_L_8, TX_L_8:  std_logic_vector (31 downto 0);
	signal credit_counter_out_8:  std_logic_vector (1 downto 0);
	signal credit_out_L_8, credit_in_L_8, valid_in_L_8, valid_out_L_8: std_logic;
	signal RX_L_9, TX_L_9:  std_logic_vector (31 downto 0);
	signal credit_counter_out_9:  std_logic_vector (1 downto 0);
	signal credit_out_L_9, credit_in_L_9, valid_in_L_9, valid_out_L_9: std_logic;
	signal RX_L_10, TX_L_10:  std_logic_vector (31 downto 0);
	signal credit_counter_out_10:  std_logic_vector (1 downto 0);
	signal credit_out_L_10, credit_in_L_10, valid_in_L_10, valid_out_L_10: std_logic;
	signal RX_L_11, TX_L_11:  std_logic_vector (31 downto 0);
	signal credit_counter_out_11:  std_logic_vector (1 downto 0);
	signal credit_out_L_11, credit_in_L_11, valid_in_L_11, valid_out_L_11: std_logic;
	signal RX_L_12, TX_L_12:  std_logic_vector (31 downto 0);
	signal credit_counter_out_12:  std_logic_vector (1 downto 0);
	signal credit_out_L_12, credit_in_L_12, valid_in_L_12, valid_out_L_12: std_logic;
	signal RX_L_13, TX_L_13:  std_logic_vector (31 downto 0);
	signal credit_counter_out_13:  std_logic_vector (1 downto 0);
	signal credit_out_L_13, credit_in_L_13, valid_in_L_13, valid_out_L_13: std_logic;
	signal RX_L_14, TX_L_14:  std_logic_vector (31 downto 0);
	signal credit_counter_out_14:  std_logic_vector (1 downto 0);
	signal credit_out_L_14, credit_in_L_14, valid_in_L_14, valid_out_L_14: std_logic;
	signal RX_L_15, TX_L_15:  std_logic_vector (31 downto 0);
	signal credit_counter_out_15:  std_logic_vector (1 downto 0);
	signal credit_out_L_15, credit_in_L_15, valid_in_L_15, valid_out_L_15: std_logic;
	--------------
	constant clk_period : time := 10 ns;
	signal reset, not_reset, clk: std_logic :='0';

	signal link_faults_0 : std_logic_vector(4 downto 0);
	signal turn_faults_0 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_0 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_0 : std_logic_vector(3 downto 0):= "1010";
	signal Reconfig_command_0 : std_logic := '0';
	signal link_faults_async_0 : std_logic_vector(4 downto 0);
	signal turn_faults_async_0 : std_logic_vector(19 downto 0);

	signal link_faults_1 : std_logic_vector(4 downto 0);
	signal turn_faults_1 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_1 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_1 : std_logic_vector(3 downto 0):= "1110";
	signal Reconfig_command_1 : std_logic := '0';
	signal link_faults_async_1 : std_logic_vector(4 downto 0);
	signal turn_faults_async_1 : std_logic_vector(19 downto 0);

	signal link_faults_2 : std_logic_vector(4 downto 0);
	signal turn_faults_2 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_2 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_2 : std_logic_vector(3 downto 0):= "1110";
	signal Reconfig_command_2 : std_logic := '0';
	signal link_faults_async_2 : std_logic_vector(4 downto 0);
	signal turn_faults_async_2 : std_logic_vector(19 downto 0);

	signal link_faults_3 : std_logic_vector(4 downto 0);
	signal turn_faults_3 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_3 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_3 : std_logic_vector(3 downto 0):= "1100";
	signal Reconfig_command_3 : std_logic := '0';
	signal link_faults_async_3 : std_logic_vector(4 downto 0);
	signal turn_faults_async_3 : std_logic_vector(19 downto 0);

	signal link_faults_4 : std_logic_vector(4 downto 0);
	signal turn_faults_4 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_4 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_4 : std_logic_vector(3 downto 0):= "1011";
	signal Reconfig_command_4 : std_logic := '0';
	signal link_faults_async_4 : std_logic_vector(4 downto 0);
	signal turn_faults_async_4 : std_logic_vector(19 downto 0);

	signal link_faults_5 : std_logic_vector(4 downto 0);
	signal turn_faults_5 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_5 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_5 : std_logic_vector(3 downto 0):= "1111";
	signal Reconfig_command_5 : std_logic := '0';
	signal link_faults_async_5 : std_logic_vector(4 downto 0);
	signal turn_faults_async_5 : std_logic_vector(19 downto 0);

	signal link_faults_6 : std_logic_vector(4 downto 0);
	signal turn_faults_6 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_6 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_6 : std_logic_vector(3 downto 0):= "1111";
	signal Reconfig_command_6 : std_logic := '0';
	signal link_faults_async_6 : std_logic_vector(4 downto 0);
	signal turn_faults_async_6 : std_logic_vector(19 downto 0);

	signal link_faults_7 : std_logic_vector(4 downto 0);
	signal turn_faults_7 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_7 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_7 : std_logic_vector(3 downto 0):= "1101";
	signal Reconfig_command_7 : std_logic := '0';
	signal link_faults_async_7 : std_logic_vector(4 downto 0);
	signal turn_faults_async_7 : std_logic_vector(19 downto 0);

	signal link_faults_8 : std_logic_vector(4 downto 0);
	signal turn_faults_8 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_8 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_8 : std_logic_vector(3 downto 0):= "1011";
	signal Reconfig_command_8 : std_logic := '0';
	signal link_faults_async_8 : std_logic_vector(4 downto 0);
	signal turn_faults_async_8 : std_logic_vector(19 downto 0);

	signal link_faults_9 : std_logic_vector(4 downto 0);
	signal turn_faults_9 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_9 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_9 : std_logic_vector(3 downto 0):= "1111";
	signal Reconfig_command_9 : std_logic := '0';
	signal link_faults_async_9 : std_logic_vector(4 downto 0);
	signal turn_faults_async_9 : std_logic_vector(19 downto 0);

	signal link_faults_10 : std_logic_vector(4 downto 0);
	signal turn_faults_10 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_10 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_10 : std_logic_vector(3 downto 0):= "1111";
	signal Reconfig_command_10 : std_logic := '0';
	signal link_faults_async_10 : std_logic_vector(4 downto 0);
	signal turn_faults_async_10 : std_logic_vector(19 downto 0);

	signal link_faults_11 : std_logic_vector(4 downto 0);
	signal turn_faults_11 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_11 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_11 : std_logic_vector(3 downto 0):= "1101";
	signal Reconfig_command_11 : std_logic := '0';
	signal link_faults_async_11 : std_logic_vector(4 downto 0);
	signal turn_faults_async_11 : std_logic_vector(19 downto 0);

	signal link_faults_12 : std_logic_vector(4 downto 0);
	signal turn_faults_12 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_12 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_12 : std_logic_vector(3 downto 0):= "0011";
	signal Reconfig_command_12 : std_logic := '0';
	signal link_faults_async_12 : std_logic_vector(4 downto 0);
	signal turn_faults_async_12 : std_logic_vector(19 downto 0);

	signal link_faults_13 : std_logic_vector(4 downto 0);
	signal turn_faults_13 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_13 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_13 : std_logic_vector(3 downto 0):= "0111";
	signal Reconfig_command_13 : std_logic := '0';
	signal link_faults_async_13 : std_logic_vector(4 downto 0);
	signal turn_faults_async_13 : std_logic_vector(19 downto 0);

	signal link_faults_14 : std_logic_vector(4 downto 0);
	signal turn_faults_14 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_14 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_14 : std_logic_vector(3 downto 0):= "0111";
	signal Reconfig_command_14 : std_logic := '0';
	signal link_faults_async_14 : std_logic_vector(4 downto 0);
	signal turn_faults_async_14 : std_logic_vector(19 downto 0);

	signal link_faults_15 : std_logic_vector(4 downto 0);
	signal turn_faults_15 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_15 : std_logic_vector(7 downto 0):= "00111100";
	signal Cx_reconf_PE_15 : std_logic_vector(3 downto 0):= "0101";
	signal Reconfig_command_15 : std_logic := '0';
	signal link_faults_async_15 : std_logic_vector(4 downto 0);
	signal turn_faults_async_15 : std_logic_vector(19 downto 0);

	-- for bubble
    signal hold_in_N_0_sig, hold_in_E_0_sig, hold_in_S_0_sig, hold_in_W_0_sig, hold_in_L_0_sig: std_logic := '1';
    signal hold_out_N_0_sig, hold_out_E_0_sig, hold_out_S_0_sig, hold_out_W_0_sig, hold_out_L_0_sig: std_logic;
    signal hold_in_N_1_sig, hold_in_E_1_sig, hold_in_S_1_sig, hold_in_W_1_sig, hold_in_L_1_sig: std_logic := '1';
    signal hold_out_N_1_sig, hold_out_E_1_sig, hold_out_S_1_sig, hold_out_W_1_sig, hold_out_L_1_sig: std_logic;
    signal hold_in_N_2_sig, hold_in_E_2_sig, hold_in_S_2_sig, hold_in_W_2_sig, hold_in_L_2_sig: std_logic := '1';
    signal hold_out_N_2_sig, hold_out_E_2_sig, hold_out_S_2_sig, hold_out_W_2_sig, hold_out_L_2_sig: std_logic;
    signal hold_in_N_3_sig, hold_in_E_3_sig, hold_in_S_3_sig, hold_in_W_3_sig, hold_in_L_3_sig: std_logic := '1';
    signal hold_out_N_3_sig, hold_out_E_3_sig, hold_out_S_3_sig, hold_out_W_3_sig, hold_out_L_3_sig: std_logic;
    signal hold_in_N_4_sig, hold_in_E_4_sig, hold_in_S_4_sig, hold_in_W_4_sig, hold_in_L_4_sig: std_logic := '1';
    signal hold_out_N_4_sig, hold_out_E_4_sig, hold_out_S_4_sig, hold_out_W_4_sig, hold_out_L_4_sig: std_logic;
    signal hold_in_N_5_sig, hold_in_E_5_sig, hold_in_S_5_sig, hold_in_W_5_sig, hold_in_L_5_sig: std_logic := '1';
    signal hold_out_N_5_sig, hold_out_E_5_sig, hold_out_S_5_sig, hold_out_W_5_sig, hold_out_L_5_sig: std_logic;
    signal hold_in_N_6_sig, hold_in_E_6_sig, hold_in_S_6_sig, hold_in_W_6_sig, hold_in_L_6_sig: std_logic := '1';
    signal hold_out_N_6_sig, hold_out_E_6_sig, hold_out_S_6_sig, hold_out_W_6_sig, hold_out_L_6_sig: std_logic;
    signal hold_in_N_7_sig, hold_in_E_7_sig, hold_in_S_7_sig, hold_in_W_7_sig, hold_in_L_7_sig: std_logic := '1';
    signal hold_out_N_7_sig, hold_out_E_7_sig, hold_out_S_7_sig, hold_out_W_7_sig, hold_out_L_7_sig: std_logic;
    signal hold_in_N_8_sig, hold_in_E_8_sig, hold_in_S_8_sig, hold_in_W_8_sig, hold_in_L_8_sig: std_logic := '1';
    signal hold_out_N_8_sig, hold_out_E_8_sig, hold_out_S_8_sig, hold_out_W_8_sig, hold_out_L_8_sig: std_logic;
    signal hold_in_N_9_sig, hold_in_E_9_sig, hold_in_S_9_sig, hold_in_W_9_sig, hold_in_L_9_sig: std_logic := '1';
    signal hold_out_N_9_sig, hold_out_E_9_sig, hold_out_S_9_sig, hold_out_W_9_sig, hold_out_L_9_sig: std_logic;
    signal hold_in_N_10_sig, hold_in_E_10_sig, hold_in_S_10_sig, hold_in_W_10_sig, hold_in_L_10_sig: std_logic := '1';
    signal hold_out_N_10_sig, hold_out_E_10_sig, hold_out_S_10_sig, hold_out_W_10_sig, hold_out_L_10_sig: std_logic;
    signal hold_in_N_11_sig, hold_in_E_11_sig, hold_in_S_11_sig, hold_in_W_11_sig, hold_in_L_11_sig: std_logic := '1';
    signal hold_out_N_11_sig, hold_out_E_11_sig, hold_out_S_11_sig, hold_out_W_11_sig, hold_out_L_11_sig: std_logic;
    signal hold_in_N_12_sig, hold_in_E_12_sig, hold_in_S_12_sig, hold_in_W_12_sig, hold_in_L_12_sig: std_logic := '1';
    signal hold_out_N_12_sig, hold_out_E_12_sig, hold_out_S_12_sig, hold_out_W_12_sig, hold_out_L_12_sig: std_logic;
    signal hold_in_N_13_sig, hold_in_E_13_sig, hold_in_S_13_sig, hold_in_W_13_sig, hold_in_L_13_sig: std_logic := '1';
    signal hold_out_N_13_sig, hold_out_E_13_sig, hold_out_S_13_sig, hold_out_W_13_sig, hold_out_L_13_sig: std_logic;
    signal hold_in_N_14_sig, hold_in_E_14_sig, hold_in_S_14_sig, hold_in_W_14_sig, hold_in_L_14_sig: std_logic := '1';
    signal hold_out_N_14_sig, hold_out_E_14_sig, hold_out_S_14_sig, hold_out_W_14_sig, hold_out_L_14_sig: std_logic;
    signal hold_in_N_15_sig, hold_in_E_15_sig, hold_in_S_15_sig, hold_in_W_15_sig, hold_in_L_15_sig: std_logic := '1';
    signal hold_out_N_15_sig, hold_out_E_15_sig, hold_out_S_15_sig, hold_out_W_15_sig, hold_out_L_15_sig: std_logic;

begin

   clk_process :process
   begin
        clk <= '0';
        wait for clk_period/2;   
        clk <= '1';
        wait for clk_period/2; 
   end process;

reset <= '1' after 1 ns;

-- instantiating the network
NoC: network_4x4 generic map (DATA_WIDTH  => 32, DATA_WIDTH_LV => 11)
port map (reset, clk, 
	RX_L_0, credit_out_L_0, valid_out_L_0, credit_in_L_0, valid_in_L_0,  TX_L_0, 
	RX_L_1, credit_out_L_1, valid_out_L_1, credit_in_L_1, valid_in_L_1,  TX_L_1, 
	RX_L_2, credit_out_L_2, valid_out_L_2, credit_in_L_2, valid_in_L_2,  TX_L_2, 
	RX_L_3, credit_out_L_3, valid_out_L_3, credit_in_L_3, valid_in_L_3,  TX_L_3, 
	RX_L_4, credit_out_L_4, valid_out_L_4, credit_in_L_4, valid_in_L_4,  TX_L_4, 
	RX_L_5, credit_out_L_5, valid_out_L_5, credit_in_L_5, valid_in_L_5,  TX_L_5, 
	RX_L_6, credit_out_L_6, valid_out_L_6, credit_in_L_6, valid_in_L_6,  TX_L_6, 
	RX_L_7, credit_out_L_7, valid_out_L_7, credit_in_L_7, valid_in_L_7,  TX_L_7, 
	RX_L_8, credit_out_L_8, valid_out_L_8, credit_in_L_8, valid_in_L_8,  TX_L_8, 
	RX_L_9, credit_out_L_9, valid_out_L_9, credit_in_L_9, valid_in_L_9,  TX_L_9, 
	RX_L_10, credit_out_L_10, valid_out_L_10, credit_in_L_10, valid_in_L_10,  TX_L_10, 
	RX_L_11, credit_out_L_11, valid_out_L_11, credit_in_L_11, valid_in_L_11,  TX_L_11, 
	RX_L_12, credit_out_L_12, valid_out_L_12, credit_in_L_12, valid_in_L_12,  TX_L_12, 
	RX_L_13, credit_out_L_13, valid_out_L_13, credit_in_L_13, valid_in_L_13,  TX_L_13, 
	RX_L_14, credit_out_L_14, valid_out_L_14, credit_in_L_14, valid_in_L_14,  TX_L_14, 
	RX_L_15, credit_out_L_15, valid_out_L_15, credit_in_L_15, valid_in_L_15,  TX_L_15, 

	link_faults_0, turn_faults_0,	Rxy_reconf_PE_0, Cx_reconf_PE_0, Reconfig_command_0, link_faults_async_0, turn_faults_async_0, 
	link_faults_1, turn_faults_1,	Rxy_reconf_PE_1, Cx_reconf_PE_1, Reconfig_command_1, link_faults_async_1, turn_faults_async_1, 
	link_faults_2, turn_faults_2,	Rxy_reconf_PE_2, Cx_reconf_PE_2, Reconfig_command_2, link_faults_async_2, turn_faults_async_2, 
	link_faults_3, turn_faults_3,	Rxy_reconf_PE_3, Cx_reconf_PE_3, Reconfig_command_3, link_faults_async_3, turn_faults_async_3, 
	link_faults_4, turn_faults_4,	Rxy_reconf_PE_4, Cx_reconf_PE_4, Reconfig_command_4, link_faults_async_4, turn_faults_async_4, 
	link_faults_5, turn_faults_5,	Rxy_reconf_PE_5, Cx_reconf_PE_5, Reconfig_command_5, link_faults_async_5, turn_faults_async_5, 
	link_faults_6, turn_faults_6,	Rxy_reconf_PE_6, Cx_reconf_PE_6, Reconfig_command_6, link_faults_async_6, turn_faults_async_6, 
	link_faults_7, turn_faults_7,	Rxy_reconf_PE_7, Cx_reconf_PE_7, Reconfig_command_7, link_faults_async_7, turn_faults_async_7, 
	link_faults_8, turn_faults_8,	Rxy_reconf_PE_8, Cx_reconf_PE_8, Reconfig_command_8, link_faults_async_8, turn_faults_async_8, 
	link_faults_9, turn_faults_9,	Rxy_reconf_PE_9, Cx_reconf_PE_9, Reconfig_command_9, link_faults_async_9, turn_faults_async_9, 
	link_faults_10, turn_faults_10,	Rxy_reconf_PE_10, Cx_reconf_PE_10, Reconfig_command_10, link_faults_async_10, turn_faults_async_10, 
	link_faults_11, turn_faults_11,	Rxy_reconf_PE_11, Cx_reconf_PE_11, Reconfig_command_11, link_faults_async_11, turn_faults_async_11, 
	link_faults_12, turn_faults_12,	Rxy_reconf_PE_12, Cx_reconf_PE_12, Reconfig_command_12, link_faults_async_12, turn_faults_async_12, 
	link_faults_13, turn_faults_13,	Rxy_reconf_PE_13, Cx_reconf_PE_13, Reconfig_command_13, link_faults_async_13, turn_faults_async_13, 
	link_faults_14, turn_faults_14,	Rxy_reconf_PE_14, Cx_reconf_PE_14, Reconfig_command_14, link_faults_async_14, turn_faults_async_14, 
	link_faults_15, turn_faults_15,	Rxy_reconf_PE_15, Cx_reconf_PE_15, Reconfig_command_15, link_faults_async_15, turn_faults_async_15,

	-- for bubbles
	hold_in_N_0_sig, hold_in_E_0_sig, hold_in_S_0_sig, hold_in_W_0_sig, hold_in_L_0_sig,
    hold_out_N_0_sig, hold_out_E_0_sig, hold_out_S_0_sig, hold_out_W_0_sig, hold_out_L_0_sig,
    hold_in_N_1_sig, hold_in_E_1_sig, hold_in_S_1_sig, hold_in_W_1_sig, hold_in_L_1_sig,
    hold_out_N_1_sig, hold_out_E_1_sig, hold_out_S_1_sig, hold_out_W_1_sig, hold_out_L_1_sig,
    hold_in_N_2_sig, hold_in_E_2_sig, hold_in_S_2_sig, hold_in_W_2_sig, hold_in_L_2_sig,
    hold_out_N_2_sig, hold_out_E_2_sig, hold_out_S_2_sig, hold_out_W_2_sig, hold_out_L_2_sig,
    hold_in_N_3_sig, hold_in_E_3_sig, hold_in_S_3_sig, hold_in_W_3_sig, hold_in_L_3_sig,
    hold_out_N_3_sig, hold_out_E_3_sig, hold_out_S_3_sig, hold_out_W_3_sig, hold_out_L_3_sig,
    hold_in_N_4_sig, hold_in_E_4_sig, hold_in_S_4_sig, hold_in_W_4_sig, hold_in_L_4_sig,
    hold_out_N_4_sig, hold_out_E_4_sig, hold_out_S_4_sig, hold_out_W_4_sig, hold_out_L_4_sig,
    hold_in_N_5_sig, hold_in_E_5_sig, hold_in_S_5_sig, hold_in_W_5_sig, hold_in_L_5_sig,
    hold_out_N_5_sig, hold_out_E_5_sig, hold_out_S_5_sig, hold_out_W_5_sig, hold_out_L_5_sig,
    hold_in_N_6_sig, hold_in_E_6_sig, hold_in_S_6_sig, hold_in_W_6_sig, hold_in_L_6_sig,
    hold_out_N_6_sig, hold_out_E_6_sig, hold_out_S_6_sig, hold_out_W_6_sig, hold_out_L_6_sig,
    hold_in_N_7_sig, hold_in_E_7_sig, hold_in_S_7_sig, hold_in_W_7_sig, hold_in_L_7_sig,
    hold_out_N_7_sig, hold_out_E_7_sig, hold_out_S_7_sig, hold_out_W_7_sig, hold_out_L_7_sig,
    hold_in_N_8_sig, hold_in_E_8_sig, hold_in_S_8_sig, hold_in_W_8_sig, hold_in_L_8_sig,
    hold_out_N_8_sig, hold_out_E_8_sig, hold_out_S_8_sig, hold_out_W_8_sig, hold_out_L_8_sig,
    hold_in_N_9_sig, hold_in_E_9_sig, hold_in_S_9_sig, hold_in_W_9_sig, hold_in_L_9_sig,
    hold_out_N_9_sig, hold_out_E_9_sig, hold_out_S_9_sig, hold_out_W_9_sig, hold_out_L_9_sig,
    hold_in_N_10_sig, hold_in_E_10_sig, hold_in_S_10_sig, hold_in_W_10_sig, hold_in_L_10_sig,
    hold_out_N_10_sig, hold_out_E_10_sig, hold_out_S_10_sig, hold_out_W_10_sig, hold_out_L_10_sig,
    hold_in_N_11_sig, hold_in_E_11_sig, hold_in_S_11_sig, hold_in_W_11_sig, hold_in_L_11_sig,
    hold_out_N_11_sig, hold_out_E_11_sig, hold_out_S_11_sig, hold_out_W_11_sig, hold_out_L_11_sig,
    hold_in_N_12_sig, hold_in_E_12_sig, hold_in_S_12_sig, hold_in_W_12_sig, hold_in_L_12_sig,
    hold_out_N_12_sig, hold_out_E_12_sig, hold_out_S_12_sig, hold_out_W_12_sig, hold_out_L_12_sig,
    hold_in_N_13_sig, hold_in_E_13_sig, hold_in_S_13_sig, hold_in_W_13_sig, hold_in_L_13_sig,
    hold_out_N_13_sig, hold_out_E_13_sig, hold_out_S_13_sig, hold_out_W_13_sig, hold_out_L_13_sig,
    hold_in_N_14_sig, hold_in_E_14_sig, hold_in_S_14_sig, hold_in_W_14_sig, hold_in_L_14_sig,
    hold_out_N_14_sig, hold_out_E_14_sig, hold_out_S_14_sig, hold_out_W_14_sig, hold_out_L_14_sig,
    hold_in_N_15_sig, hold_in_E_15_sig, hold_in_S_15_sig, hold_in_W_15_sig, hold_in_L_15_sig,
    hold_out_N_15_sig, hold_out_E_15_sig, hold_out_S_15_sig, hold_out_W_15_sig, hold_out_L_15_sig
        ); 
not_reset <= not reset; 

-- connecting the packet generators
credit_counter_control(clk, credit_out_L_0, valid_in_L_0, credit_counter_out_0);
gen_random_packet(4, 100, 0, 45, 8, 8, 10000 ns, clk, credit_counter_out_0, valid_in_L_0, RX_L_0);

credit_counter_control(clk, credit_out_L_1, valid_in_L_1, credit_counter_out_1);
gen_random_packet(4, 100, 1, 29, 8, 8, 10000 ns, clk, credit_counter_out_1, valid_in_L_1, RX_L_1);

credit_counter_control(clk, credit_out_L_2, valid_in_L_2, credit_counter_out_2);
gen_random_packet(4, 100, 2, 34, 8, 8, 10000 ns, clk, credit_counter_out_2, valid_in_L_2, RX_L_2);

credit_counter_control(clk, credit_out_L_3, valid_in_L_3, credit_counter_out_3);
gen_random_packet(4, 100, 3, 23, 8, 8, 10000 ns, clk, credit_counter_out_3, valid_in_L_3, RX_L_3);

credit_counter_control(clk, credit_out_L_4, valid_in_L_4, credit_counter_out_4);
gen_random_packet(4, 100, 4, 5, 8, 8, 10000 ns, clk, credit_counter_out_4, valid_in_L_4, RX_L_4);

credit_counter_control(clk, credit_out_L_5, valid_in_L_5, credit_counter_out_5);
gen_random_packet(4, 100, 5, 35, 8, 8, 10000 ns, clk, credit_counter_out_5, valid_in_L_5, RX_L_5);

credit_counter_control(clk, credit_out_L_6, valid_in_L_6, credit_counter_out_6);
gen_random_packet(4, 100, 6, 42, 8, 8, 10000 ns, clk, credit_counter_out_6, valid_in_L_6, RX_L_6);

credit_counter_control(clk, credit_out_L_7, valid_in_L_7, credit_counter_out_7);
gen_random_packet(4, 100, 7, 9, 8, 8, 10000 ns, clk, credit_counter_out_7, valid_in_L_7, RX_L_7);

credit_counter_control(clk, credit_out_L_8, valid_in_L_8, credit_counter_out_8);
gen_random_packet(4, 100, 8, 5, 8, 8, 10000 ns, clk, credit_counter_out_8, valid_in_L_8, RX_L_8);

credit_counter_control(clk, credit_out_L_9, valid_in_L_9, credit_counter_out_9);
gen_random_packet(4, 100, 9, 30, 8, 8, 10000 ns, clk, credit_counter_out_9, valid_in_L_9, RX_L_9);

credit_counter_control(clk, credit_out_L_10, valid_in_L_10, credit_counter_out_10);
gen_random_packet(4, 100, 10, 43, 8, 8, 10000 ns, clk, credit_counter_out_10, valid_in_L_10, RX_L_10);

credit_counter_control(clk, credit_out_L_11, valid_in_L_11, credit_counter_out_11);
gen_random_packet(4, 100, 11, 31, 8, 8, 10000 ns, clk, credit_counter_out_11, valid_in_L_11, RX_L_11);

credit_counter_control(clk, credit_out_L_12, valid_in_L_12, credit_counter_out_12);
gen_random_packet(4, 100, 12, 29, 8, 8, 10000 ns, clk, credit_counter_out_12, valid_in_L_12, RX_L_12);

credit_counter_control(clk, credit_out_L_13, valid_in_L_13, credit_counter_out_13);
gen_random_packet(4, 100, 13, 8, 8, 8, 10000 ns, clk, credit_counter_out_13, valid_in_L_13, RX_L_13);

credit_counter_control(clk, credit_out_L_14, valid_in_L_14, credit_counter_out_14);
gen_random_packet(4, 100, 14, 27, 8, 8, 10000 ns, clk, credit_counter_out_14, valid_in_L_14, RX_L_14);

credit_counter_control(clk, credit_out_L_15, valid_in_L_15, credit_counter_out_15);
gen_random_packet(4, 100, 15, 7, 8, 8, 10000 ns, clk, credit_counter_out_15, valid_in_L_15, RX_L_15);


-- connecting the packet receivers
get_packet(32, 5, 0, clk, credit_in_L_0, valid_out_L_0,  TX_L_0);
get_packet(32, 5, 1, clk, credit_in_L_1, valid_out_L_1,  TX_L_1);
get_packet(32, 5, 2, clk, credit_in_L_2, valid_out_L_2,  TX_L_2);
get_packet(32, 5, 3, clk, credit_in_L_3, valid_out_L_3,  TX_L_3);
get_packet(32, 5, 4, clk, credit_in_L_4, valid_out_L_4,  TX_L_4);
get_packet(32, 5, 5, clk, credit_in_L_5, valid_out_L_5,  TX_L_5);
get_packet(32, 5, 6, clk, credit_in_L_6, valid_out_L_6,  TX_L_6);
get_packet(32, 5, 7, clk, credit_in_L_7, valid_out_L_7,  TX_L_7);
get_packet(32, 5, 8, clk, credit_in_L_8, valid_out_L_8,  TX_L_8);
get_packet(32, 5, 9, clk, credit_in_L_9, valid_out_L_9,  TX_L_9);
get_packet(32, 5, 10, clk, credit_in_L_10, valid_out_L_10,  TX_L_10);
get_packet(32, 5, 11, clk, credit_in_L_11, valid_out_L_11,  TX_L_11);
get_packet(32, 5, 12, clk, credit_in_L_12, valid_out_L_12,  TX_L_12);
get_packet(32, 5, 13, clk, credit_in_L_13, valid_out_L_13,  TX_L_13);
get_packet(32, 5, 14, clk, credit_in_L_14, valid_out_L_14,  TX_L_14);
get_packet(32, 5, 15, clk, credit_in_L_15, valid_out_L_15,  TX_L_15);


end;
